`timescale 1ns / 1ps

module OR(
	   input [31:0] I1,
	   input [31:0] I2,
	   output [31:0] O);
              	   
assign O = I1 | I2;
endmodule